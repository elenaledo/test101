a<= b
