Elena says "duck you", and TuanPham feels painful :)
