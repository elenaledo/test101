First by Elena
