feature for test
