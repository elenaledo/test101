A feature by Elena
