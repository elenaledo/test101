Elena create mem :)
