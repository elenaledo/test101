Elena says "duck you", and TuanPham feels painful :)
Elena says "Marcus has 9 inch", and TuanPham feels emotional damage :)
