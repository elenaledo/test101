First by Elena
Second by Elena
