Elena is stoopid
