Rio is not stoopid but just retard
